/* Environment class will instantiate and connect generator, driver, monitor , scoreboard.
It will also manage all the mailbox 