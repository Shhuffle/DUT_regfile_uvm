/* What an Environment Class Does:
1. Instantiates components: generator, driver, monitor, scoreboard
2. Creates and shares common resources (like mailbox, virtual interface)
3. Starts the run methods of these components
4. Acts as a container to manage the testbench flow*/



